LPFILTER.CIR - SIMPLE RC LOW-PASS FILTER
VS	1	0	AC	1	SIN(0VOFF 1VPEAK   2KHZ)
R1	1	2	1K
C1	2	0	0.032UF
*
* ANALYSIS
.AC 	DEC 	5 10 10MEG
.TRAN 	5US  500US
* VIEW RESULTS
.PRINT	AC 	VM(2) VP(2)
.PLOT	AC	VM(2) VP(2)
.PRINT	TRAN 	V(1) V(2)
.PLOT	TRAN 	V(1) V(2)
.PROBE
.END
